module Checkkeypad(clk,rst,keypadRow,keypadCol,keypadBuf);

input clk,rst;
input [3:0] keypadCol;
output [3:0] keypadRow;
output [3:0] keypadBuf;

reg [3:0] keypadRow;
reg [3:0] keypadBuf;
reg [31:0] keypadDelay;

always@(posedge clk or negedge rst)
begin
   if(!rst)
	begin
	   keypadRow<=4'b1110;
		keypadBuf<=4'b0000;
		keypadDelay<=31'd0;
	end
	else
	begin
	   //if(keypadDelay==`TimeExpire_KEY)
		begin
		   keypadDelay=31'd0;
			case({keypadRow,keypadCol})
			   8'b1110_1110:keypadBuf<=4'h7;
				8'b1110_1101:keypadBuf<=4'h4;
				8'b1110_1011:keypadBuf<=4'h1;
				8'b1110_0111:keypadBuf<=4'h0;
				8'b1101_1110:keypadBuf<=4'h8;
				8'b1101_1101:keypadBuf<=4'h5;
				8'b1101_1011:keypadBuf<=4'h2;
				8'b1101_0111:keypadBuf<=4'ha;
				8'b1011_1110:keypadBuf<=4'h9;
				8'b1011_1101:keypadBuf<=4'h6;
				8'b1011_1011:keypadBuf<=4'h3;
				8'b1011_0111:keypadBuf<=4'hb;
				8'b0111_1110:keypadBuf<=4'hc;
				8'b0111_1101:keypadBuf<=4'hd;
				8'b0111_1011:keypadBuf<=4'he;
				8'b0111_0111:keypadBuf<=4'hf;
				default     :keypadBuf<=keypadBuf;
			endcase
		case(keypadRow)
		   4'b1110:keypadRow<=4'b1101;
			4'b1101:keypadRow<=4'b1011;
			4'b1011:keypadRow<=4'b0111;
			4'b0111:keypadRow<=4'b1110;
			default:keypadRow<=4'b1110;
		endcase
	   end
	//else
	  // keypadDelay<=keypadDelay+1'b1;
	end
end
endmodule 